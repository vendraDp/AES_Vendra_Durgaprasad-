module Mod1 (Sin, Sout);

input  [0:7] Sin;
output [0:7] Sout;

assign Sout[0:7] = Sin[0:7];

endmodule
